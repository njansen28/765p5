module lfsr247(clk, bist_en, rst_l, value);
	input clk, bist_en, rst_l;
	output [246:0] value;

  // init stuff
  //wire s0_l;// set to zero, asserted low
  //not g0 (s0_l, init);

  // tap stuff
  wire tapping165, bist_clk, init_bist, init_state, n_init_state, init;
  xor g1 (tapping165, value[0], value[165]);
  and bist_clk_and(bist_clk, clk, bist_en);
  
  //stuff to init only at start
  dff_r bist_init_ff(init_state, clk, rst_l, bist_en);
  not bistn(n_init_state, init_state);
  and bist_init_and(init, n_init_state, bist_en);
  not initn(init_bist, init);
  // dff stuff

  dff0 d000 (value[  0], bist_clk, value[  1], init_bist);
  dff1 d001 (value[  1], bist_clk, value[  2], init_bist);
  dff1 d002 (value[  2], bist_clk, value[  3], init_bist);
  dff1 d003 (value[  3], bist_clk, value[  4], init_bist);
  dff0 d004 (value[  4], bist_clk, value[  5], init_bist);
  dff0 d005 (value[  5], bist_clk, value[  6], init_bist);
  dff0 d006 (value[  6], bist_clk, value[  7], init_bist);
  dff0 d007 (value[  7], bist_clk, value[  8], init_bist);
  dff0 d008 (value[  8], bist_clk, value[  9], init_bist);
  dff1 d009 (value[  9], bist_clk, value[ 10], init_bist);
                                        
  dff0 d010 (value[ 10], bist_clk, value[ 11], init_bist);
  dff0 d011 (value[ 11], bist_clk, value[ 12], init_bist);
  dff1 d012 (value[ 12], bist_clk, value[ 13], init_bist);
  dff0 d013 (value[ 13], bist_clk, value[ 14], init_bist);
  dff1 d014 (value[ 14], bist_clk, value[ 15], init_bist);
  dff0 d015 (value[ 15], bist_clk, value[ 16], init_bist);
  dff1 d016 (value[ 16], bist_clk, value[ 17], init_bist);
  dff0 d017 (value[ 17], bist_clk, value[ 18], init_bist);
  dff1 d018 (value[ 18], bist_clk, value[ 19], init_bist);
  dff1 d019 (value[ 19], bist_clk, value[ 20], init_bist);
                                        
  dff0 d020 (value[ 20], bist_clk, value[ 21], init_bist);
  dff1 d021 (value[ 21], bist_clk, value[ 22], init_bist);
  dff0 d022 (value[ 22], bist_clk, value[ 23], init_bist);
  dff0 d023 (value[ 23], bist_clk, value[ 24], init_bist);
  dff1 d024 (value[ 24], bist_clk, value[ 25], init_bist);
  dff0 d025 (value[ 25], bist_clk, value[ 26], init_bist);
  dff0 d026 (value[ 26], bist_clk, value[ 27], init_bist);
  dff0 d027 (value[ 27], bist_clk, value[ 28], init_bist);
  dff0 d028 (value[ 28], bist_clk, value[ 29], init_bist);
  dff1 d029 (value[ 29], bist_clk, value[ 30], init_bist);
                                        
  dff1 d030 (value[ 30], bist_clk, value[ 31], init_bist);
  dff0 d031 (value[ 31], bist_clk, value[ 32], init_bist);
  dff0 d032 (value[ 32], bist_clk, value[ 33], init_bist);
  dff0 d033 (value[ 33], bist_clk, value[ 34], init_bist);
  dff1 d034 (value[ 34], bist_clk, value[ 35], init_bist);
  dff1 d035 (value[ 35], bist_clk, value[ 36], init_bist);
  dff1 d036 (value[ 36], bist_clk, value[ 37], init_bist);
  dff0 d037 (value[ 37], bist_clk, value[ 38], init_bist);
  dff1 d038 (value[ 38], bist_clk, value[ 39], init_bist);
  dff0 d039 (value[ 39], bist_clk, value[ 40], init_bist);
                                        
  dff0 d040 (value[ 40], bist_clk, value[ 41], init_bist);
  dff0 d041 (value[ 41], bist_clk, value[ 42], init_bist);
  dff1 d042 (value[ 42], bist_clk, value[ 43], init_bist);
  dff0 d043 (value[ 43], bist_clk, value[ 44], init_bist);
  dff1 d044 (value[ 44], bist_clk, value[ 45], init_bist);
  dff1 d045 (value[ 45], bist_clk, value[ 46], init_bist);
  dff0 d046 (value[ 46], bist_clk, value[ 47], init_bist);
  dff0 d047 (value[ 47], bist_clk, value[ 48], init_bist);
  dff0 d048 (value[ 48], bist_clk, value[ 49], init_bist);
  dff0 d049 (value[ 49], bist_clk, value[ 50], init_bist);
                                        
  dff0 d050 (value[ 50], bist_clk, value[ 51], init_bist);
  dff1 d051 (value[ 51], bist_clk, value[ 52], init_bist);
  dff0 d052 (value[ 52], bist_clk, value[ 53], init_bist);
  dff1 d053 (value[ 53], bist_clk, value[ 54], init_bist);
  dff1 d054 (value[ 54], bist_clk, value[ 55], init_bist);
  dff1 d055 (value[ 55], bist_clk, value[ 56], init_bist);
  dff1 d056 (value[ 56], bist_clk, value[ 57], init_bist);
  dff1 d057 (value[ 57], bist_clk, value[ 58], init_bist);
  dff1 d058 (value[ 58], bist_clk, value[ 59], init_bist);
  dff1 d059 (value[ 59], bist_clk, value[ 60], init_bist);
                                        
  dff0 d060 (value[ 60], bist_clk, value[ 61], init_bist);
  dff0 d061 (value[ 61], bist_clk, value[ 62], init_bist);
  dff1 d062 (value[ 62], bist_clk, value[ 63], init_bist);
  dff1 d063 (value[ 63], bist_clk, value[ 64], init_bist);
  dff1 d064 (value[ 64], bist_clk, value[ 65], init_bist);
  dff1 d065 (value[ 65], bist_clk, value[ 66], init_bist);
  dff1 d066 (value[ 66], bist_clk, value[ 67], init_bist);
  dff1 d067 (value[ 67], bist_clk, value[ 68], init_bist);
  dff1 d068 (value[ 68], bist_clk, value[ 69], init_bist);
  dff0 d069 (value[ 69], bist_clk, value[ 70], init_bist);
                                        
  dff1 d070 (value[ 70], bist_clk, value[ 71], init_bist);
  dff0 d071 (value[ 71], bist_clk, value[ 72], init_bist);
  dff0 d072 (value[ 72], bist_clk, value[ 73], init_bist);
  dff1 d073 (value[ 73], bist_clk, value[ 74], init_bist);
  dff0 d074 (value[ 74], bist_clk, value[ 75], init_bist);
  dff1 d075 (value[ 75], bist_clk, value[ 76], init_bist);
  dff1 d076 (value[ 76], bist_clk, value[ 77], init_bist);
  dff0 d077 (value[ 77], bist_clk, value[ 78], init_bist);
  dff1 d078 (value[ 78], bist_clk, value[ 79], init_bist);
  dff0 d079 (value[ 79], bist_clk, value[ 80], init_bist);
                                        
  dff0 d080 (value[ 80], bist_clk, value[ 81], init_bist);
  dff0 d081 (value[ 81], bist_clk, value[ 82], init_bist);
  dff0 d082 (value[ 82], bist_clk, value[ 83], init_bist);
  dff0 d083 (value[ 83], bist_clk, value[ 84], init_bist);
  dff0 d084 (value[ 84], bist_clk, value[ 85], init_bist);
  dff1 d085 (value[ 85], bist_clk, value[ 86], init_bist);
  dff0 d086 (value[ 86], bist_clk, value[ 87], init_bist);
  dff1 d087 (value[ 87], bist_clk, value[ 88], init_bist);
  dff0 d088 (value[ 88], bist_clk, value[ 89], init_bist);
  dff0 d089 (value[ 89], bist_clk, value[ 90], init_bist);
                                        
  dff1 d090 (value[ 90], bist_clk, value[ 91], init_bist);
  dff1 d091 (value[ 91], bist_clk, value[ 92], init_bist);
  dff1 d092 (value[ 92], bist_clk, value[ 93], init_bist);
  dff1 d093 (value[ 93], bist_clk, value[ 94], init_bist);
  dff1 d094 (value[ 94], bist_clk, value[ 95], init_bist);
  dff0 d095 (value[ 95], bist_clk, value[ 96], init_bist);
  dff0 d096 (value[ 96], bist_clk, value[ 97], init_bist);
  dff0 d097 (value[ 97], bist_clk, value[ 98], init_bist);
  dff0 d098 (value[ 98], bist_clk, value[ 99], init_bist);
  dff0 d099 (value[ 99], bist_clk, value[100], init_bist);
                                         
                                        
  dff0 d100 (value[100], bist_clk, value[101], init_bist);
  dff0 d101 (value[101], bist_clk, value[102], init_bist);
  dff0 d102 (value[102], bist_clk, value[103], init_bist);
  dff0 d103 (value[103], bist_clk, value[104], init_bist);
  dff1 d104 (value[104], bist_clk, value[105], init_bist);
  dff1 d105 (value[105], bist_clk, value[106], init_bist);
  dff0 d106 (value[106], bist_clk, value[107], init_bist);
  dff1 d107 (value[107], bist_clk, value[108], init_bist);
  dff0 d108 (value[108], bist_clk, value[109], init_bist);
  dff1 d109 (value[109], bist_clk, value[110], init_bist);
                                        
  dff1 d110 (value[110], bist_clk, value[111], init_bist);
  dff1 d111 (value[111], bist_clk, value[112], init_bist);
  dff1 d112 (value[112], bist_clk, value[113], init_bist);
  dff1 d113 (value[113], bist_clk, value[114], init_bist);
  dff1 d114 (value[114], bist_clk, value[115], init_bist);
  dff1 d115 (value[115], bist_clk, value[116], init_bist);
  dff1 d116 (value[116], bist_clk, value[117], init_bist);
  dff1 d117 (value[117], bist_clk, value[118], init_bist);
  dff0 d118 (value[118], bist_clk, value[119], init_bist);
  dff1 d119 (value[119], bist_clk, value[120], init_bist);
                                       
  dff0 d120 (value[120], bist_clk, value[121], init_bist);
  dff0 d121 (value[121], bist_clk, value[122], init_bist);
  dff0 d122 (value[122], bist_clk, value[123], init_bist);
  dff0 d123 (value[123], bist_clk, value[124], init_bist);
  dff0 d124 (value[124], bist_clk, value[125], init_bist);
  dff0 d125 (value[125], bist_clk, value[126], init_bist);
  dff1 d126 (value[126], bist_clk, value[127], init_bist);
  dff0 d127 (value[127], bist_clk, value[128], init_bist);
  dff0 d128 (value[128], bist_clk, value[129], init_bist);
  dff1 d129 (value[129], bist_clk, value[130], init_bist);
                                        
  dff1 d130 (value[130], bist_clk, value[131], init_bist);
  dff1 d131 (value[131], bist_clk, value[132], init_bist);
  dff0 d132 (value[132], bist_clk, value[133], init_bist);
  dff1 d133 (value[133], bist_clk, value[134], init_bist);
  dff0 d134 (value[134], bist_clk, value[135], init_bist);
  dff1 d135 (value[135], bist_clk, value[136], init_bist);
  dff1 d136 (value[136], bist_clk, value[137], init_bist);
  dff0 d137 (value[137], bist_clk, value[138], init_bist);
  dff1 d138 (value[138], bist_clk, value[139], init_bist);
  dff0 d139 (value[139], bist_clk, value[140], init_bist);
                                        
  dff1 d140 (value[140], bist_clk, value[141], init_bist);
  dff0 d141 (value[141], bist_clk, value[142], init_bist);
  dff1 d142 (value[142], bist_clk, value[143], init_bist);
  dff1 d143 (value[143], bist_clk, value[144], init_bist);
  dff1 d144 (value[144], bist_clk, value[145], init_bist);
  dff1 d145 (value[145], bist_clk, value[146], init_bist);
  dff1 d146 (value[146], bist_clk, value[147], init_bist);
  dff0 d147 (value[147], bist_clk, value[148], init_bist);
  dff1 d148 (value[148], bist_clk, value[149], init_bist);
  dff0 d149 (value[149], bist_clk, value[150], init_bist);
                                        
  dff1 d150 (value[150], bist_clk, value[151], init_bist);
  dff0 d151 (value[151], bist_clk, value[152], init_bist);
  dff1 d152 (value[152], bist_clk, value[153], init_bist);
  dff0 d153 (value[153], bist_clk, value[154], init_bist);
  dff1 d154 (value[154], bist_clk, value[155], init_bist);
  dff1 d155 (value[155], bist_clk, value[156], init_bist);
  dff0 d156 (value[156], bist_clk, value[157], init_bist);
  dff0 d157 (value[157], bist_clk, value[158], init_bist);
  dff0 d158 (value[158], bist_clk, value[159], init_bist);
  dff0 d159 (value[159], bist_clk, value[160], init_bist);
                                        
  dff1 d160 (value[160], bist_clk, value[161], init_bist);
  dff0 d161 (value[161], bist_clk, value[162], init_bist);
  dff1 d162 (value[162], bist_clk, value[163], init_bist);
  dff1 d163 (value[163], bist_clk, value[164], init_bist);
  dff1 d164 (value[164], bist_clk, tapping165, init_bist); // tap 165
  dff0 d165 (value[165], bist_clk, value[166], init_bist);
  dff1 d166 (value[166], bist_clk, value[167], init_bist);
  dff1 d167 (value[167], bist_clk, value[168], init_bist);
  dff0 d168 (value[168], bist_clk, value[169], init_bist);
  dff1 d169 (value[169], bist_clk, value[170], init_bist);
                                        
  dff0 d170 (value[170], bist_clk, value[171], init_bist);
  dff1 d171 (value[171], bist_clk, value[172], init_bist);
  dff1 d172 (value[172], bist_clk, value[173], init_bist);
  dff1 d173 (value[173], bist_clk, value[174], init_bist);
  dff1 d174 (value[174], bist_clk, value[175], init_bist);
  dff0 d175 (value[175], bist_clk, value[176], init_bist);
  dff1 d176 (value[176], bist_clk, value[177], init_bist);
  dff1 d177 (value[177], bist_clk, value[178], init_bist);
  dff0 d178 (value[178], bist_clk, value[179], init_bist);
  dff0 d179 (value[179], bist_clk, value[180], init_bist);
                                        
  dff1 d180 (value[180], bist_clk, value[181], init_bist);
  dff0 d181 (value[181], bist_clk, value[182], init_bist);
  dff0 d182 (value[182], bist_clk, value[183], init_bist);
  dff0 d183 (value[183], bist_clk, value[184], init_bist);
  dff1 d184 (value[184], bist_clk, value[185], init_bist);
  dff1 d185 (value[185], bist_clk, value[186], init_bist);
  dff1 d186 (value[186], bist_clk, value[187], init_bist);
  dff0 d187 (value[187], bist_clk, value[188], init_bist);
  dff0 d188 (value[188], bist_clk, value[189], init_bist);
  dff1 d189 (value[189], bist_clk, value[190], init_bist);
                                         
  dff1 d190 (value[190], bist_clk, value[191], init_bist);
  dff0 d191 (value[191], bist_clk, value[192], init_bist);
  dff1 d192 (value[192], bist_clk, value[193], init_bist);
  dff0 d193 (value[193], bist_clk, value[194], init_bist);
  dff0 d194 (value[194], bist_clk, value[195], init_bist);
  dff1 d195 (value[195], bist_clk, value[196], init_bist);
  dff1 d196 (value[196], bist_clk, value[197], init_bist);
  dff0 d197 (value[197], bist_clk, value[198], init_bist);
  dff0 d198 (value[198], bist_clk, value[199], init_bist);
  dff1 d199 (value[199], bist_clk, value[200], init_bist);
                                         
                                        
  dff1 d200 (value[200], bist_clk, value[201], init_bist);
  dff0 d201 (value[201], bist_clk, value[202], init_bist);
  dff1 d202 (value[202], bist_clk, value[203], init_bist);
  dff0 d203 (value[203], bist_clk, value[204], init_bist);
  dff1 d204 (value[204], bist_clk, value[205], init_bist);
  dff1 d205 (value[205], bist_clk, value[206], init_bist);
  dff0 d206 (value[206], bist_clk, value[207], init_bist);
  dff0 d207 (value[207], bist_clk, value[208], init_bist);
  dff1 d208 (value[208], bist_clk, value[209], init_bist);
  dff1 d209 (value[209], bist_clk, value[210], init_bist);
                                        
  dff1 d210 (value[210], bist_clk, value[211], init_bist);
  dff0 d211 (value[211], bist_clk, value[212], init_bist);
  dff1 d212 (value[212], bist_clk, value[213], init_bist);
  dff1 d213 (value[213], bist_clk, value[214], init_bist);
  dff1 d214 (value[214], bist_clk, value[215], init_bist);
  dff0 d215 (value[215], bist_clk, value[216], init_bist);
  dff0 d216 (value[216], bist_clk, value[217], init_bist);
  dff1 d217 (value[217], bist_clk, value[218], init_bist);
  dff1 d218 (value[218], bist_clk, value[219], init_bist);
  dff0 d219 (value[219], bist_clk, value[220], init_bist);
                                        
  dff0 d220 (value[220], bist_clk, value[221], init_bist);
  dff1 d221 (value[221], bist_clk, value[222], init_bist);
  dff1 d222 (value[222], bist_clk, value[223], init_bist);
  dff1 d223 (value[223], bist_clk, value[224], init_bist);
  dff1 d224 (value[224], bist_clk, value[225], init_bist);
  dff0 d225 (value[225], bist_clk, value[226], init_bist);
  dff0 d226 (value[226], bist_clk, value[227], init_bist);
  dff1 d227 (value[227], bist_clk, value[228], init_bist);
  dff0 d228 (value[228], bist_clk, value[229], init_bist);
  dff1 d229 (value[229], bist_clk, value[230], init_bist);
                                        
  dff0 d230 (value[230], bist_clk, value[231], init_bist);
  dff0 d231 (value[231], bist_clk, value[232], init_bist);
  dff0 d232 (value[232], bist_clk, value[233], init_bist);
  dff0 d233 (value[233], bist_clk, value[234], init_bist);
  dff0 d234 (value[234], bist_clk, value[235], init_bist);
  dff0 d235 (value[235], bist_clk, value[236], init_bist);
  dff0 d236 (value[236], bist_clk, value[237], init_bist);
  dff1 d237 (value[237], bist_clk, value[238], init_bist);
  dff1 d238 (value[238], bist_clk, value[239], init_bist);
  dff1 d239 (value[239], bist_clk, value[240], init_bist);
                                        
  dff1 d240 (value[240], bist_clk, value[241], init_bist);
  dff0 d241 (value[241], bist_clk, value[242], init_bist);
  dff1 d242 (value[242], bist_clk, value[243], init_bist);
  dff0 d243 (value[243], bist_clk, value[244], init_bist);
  dff0 d244 (value[244], bist_clk, value[245], init_bist);
  dff1 d245 (value[245], bist_clk, value[246], init_bist);
  dff1 d246 (value[246], bist_clk, value[  0], init_bist); // tap 247 (tapping 0)
     
endmodule

`default_nettype wire
// cost 1.2
module dff0 (q, clock, data, rst_l);
  input clock, data, rst_l;
  output q;
  
  wire d;

  and (d, data, rst_l);
  dff f (q, clock, d);

endmodule

// cost 1.2
module dff1 (q, clock, data, rst_l);
  input clock, data, rst_l;
  output q;
  
  wire d, rst;
  

  not n0(rst, rst_l);  
  or(d, data, rst);
  dff f (q, clock, d);

endmodule

module xor125(
	input [124:0] x,
	output y
	);
	xor x0(y,
		x[  0],
		x[  1],
		x[  2],
		x[  3],
		x[  4],
		x[  5],
		x[  6],
		x[  7],
		x[  8],
		x[  9],
		
		x[ 10],
		x[ 11],
		x[ 12],
		x[ 13],
		x[ 14],
		x[ 15],
		x[ 16],
		x[ 17],
		x[ 18],
		x[ 19],
		
		x[ 20],
		x[ 21],
		x[ 22],
		x[ 23],
		x[ 24],
		x[ 25],
		x[ 26],
		x[ 27],
		x[ 28],
		x[ 29],
		
		x[ 30],
		x[ 31],
		x[ 32],
		x[ 33],
		x[ 34],
		x[ 35],
		x[ 36],
		x[ 37],
		x[ 38],
		x[ 39],
		
		x[ 40],
		x[ 41],
		x[ 42],
		x[ 43],
		x[ 44],
		x[ 45],
		x[ 46],
		x[ 47],
		x[ 48],
		x[ 49],
		
		x[ 50],
		x[ 51],
		x[ 52],
		x[ 53],
		x[ 54],
		x[ 55],
		x[ 56],
		x[ 57],
		x[ 58],
		x[ 59],
		
		x[ 60],
		x[ 61],
		x[ 62],
		x[ 63],
		x[ 64],
		x[ 65],
		x[ 66],
		x[ 67],
		x[ 68],
		x[ 69],
		
		x[ 70],
		x[ 71],
		x[ 72],
		x[ 73],
		x[ 74],
		x[ 75],
		x[ 76],
		x[ 77],
		x[ 78],
		x[ 79],
		
		x[ 80],
		x[ 81],
		x[ 82],
		x[ 83],
		x[ 84],
		x[ 85],
		x[ 86],
		x[ 87],
		x[ 88],
		x[ 89],
		
		x[ 90],
		x[ 91],
		x[ 92],
		x[ 93],
		x[ 94],
		x[ 95],
		x[ 96],
		x[ 97],
		x[ 98],
		x[ 99],
		
		
		x[100],
		x[101],
		x[102],
		x[103],
		x[104],
		x[105],
		x[106],
		x[107],
		x[108],
		x[109],
		
		x[110],
		x[111],
		x[112],
		x[113],
		x[114],
		x[115],
		x[116],
		x[117],
		x[118],
		x[119],
		
		x[120],
		x[121],
		x[122],
		x[123],
		x[124]);
			
	
endmodule // xor125



module xor250(
  input [249:0] x,
  output y
);

xor(
  y,

  x[  0],
  x[  1],
  x[  2],
  x[  3],
  x[  4],
  x[  5],
  x[  6],
  x[  7],
  x[  8],
  x[  9],

  x[ 10],
  x[ 11],
  x[ 12],
  x[ 13],
  x[ 14],
  x[ 15],
  x[ 16],
  x[ 17],
  x[ 18],
  x[ 19],

  x[ 20],
  x[ 21],
  x[ 22],
  x[ 23],
  x[ 24],
  x[ 25],
  x[ 26],
  x[ 27],
  x[ 28],
  x[ 29],

  x[ 30],
  x[ 31],
  x[ 32],
  x[ 33],
  x[ 34],
  x[ 35],
  x[ 36],
  x[ 37],
  x[ 38],
  x[ 39],

  x[ 40],
  x[ 41],
  x[ 42],
  x[ 43],
  x[ 44],
  x[ 45],
  x[ 46],
  x[ 47],
  x[ 48],
  x[ 49],

  x[ 50],
  x[ 51],
  x[ 52],
  x[ 53],
  x[ 54],
  x[ 55],
  x[ 56],
  x[ 57],
  x[ 58],
  x[ 59],

  x[ 60],
  x[ 61],
  x[ 62],
  x[ 63],
  x[ 64],
  x[ 65],
  x[ 66],
  x[ 67],
  x[ 68],
  x[ 69],

  x[ 70],
  x[ 71],
  x[ 72],
  x[ 73],
  x[ 74],
  x[ 75],
  x[ 76],
  x[ 77],
  x[ 78],
  x[ 79],

  x[ 80],
  x[ 81],
  x[ 82],
  x[ 83],
  x[ 84],
  x[ 85],
  x[ 86],
  x[ 87],
  x[ 88],
  x[ 89],

  x[ 90],
  x[ 91],
  x[ 92],
  x[ 93],
  x[ 94],
  x[ 95],
  x[ 96],
  x[ 97],
  x[ 98],
  x[ 99],


  x[100],
  x[101],
  x[102],
  x[103],
  x[104],
  x[105],
  x[106],
  x[107],
  x[108],
  x[109],

  x[110],
  x[111],
  x[112],
  x[113],
  x[114],
  x[115],
  x[116],
  x[117],
  x[118],
  x[119],

  x[120],
  x[121],
  x[122],
  x[123],
  x[124],
  x[125],
  x[126],
  x[127],
  x[128],
  x[129],

  x[130],
  x[131],
  x[132],
  x[133],
  x[134],
  x[135],
  x[136],
  x[137],
  x[138],
  x[139],

  x[140],
  x[141],
  x[142],
  x[143],
  x[144],
  x[145],
  x[146],
  x[147],
  x[148],
  x[149],

  x[150],
  x[151],
  x[152],
  x[153],
  x[154],
  x[155],
  x[156],
  x[157],
  x[158],
  x[159],

  x[160],
  x[161],
  x[162],
  x[163],
  x[164],
  x[165],
  x[166],
  x[167],
  x[168],
  x[169],

  x[170],
  x[171],
  x[172],
  x[173],
  x[174],
  x[175],
  x[176],
  x[177],
  x[178],
  x[179],

  x[180],
  x[181],
  x[182],
  x[183],
  x[184],
  x[185],
  x[186],
  x[187],
  x[188],
  x[189],

  x[190],
  x[191],
  x[192],
  x[193],
  x[194],
  x[195],
  x[196],
  x[197],
  x[198],
  x[199],

  x[200],
  x[201],
  x[202],
  x[203],
  x[204],
  x[205],
  x[206],
  x[207],
  x[208],
  x[209],

  x[210],
  x[211],
  x[212],
  x[213],
  x[214],
  x[215],
  x[216],
  x[217],
  x[218],
  x[219],

  x[220],
  x[221],
  x[222],
  x[223],
  x[224],
  x[225],
  x[226],
  x[227],
  x[228],
  x[229],

  x[230],
  x[231],
  x[232],
  x[233],
  x[234],
  x[235],
  x[236],
  x[237],
  x[238],
  x[239],

  x[240],
  x[241],
  x[242],
  x[243],
  x[244],
  x[245],
  x[246]
);
endmodule
